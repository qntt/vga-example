
module equal1 (
	source,
	probe);	

	output	[0:0]	source;
	input	[49:0]	probe;
endmodule
