module skeleton(resetn, 
	ps2_clock, ps2_data, 										// ps2 related I/O
	debug_data_in, debug_addr, leds, 						// extra debugging ports
	lcd_data, lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon,// LCD info
	seg1, seg2, seg3, seg4, seg5, seg6, seg7, seg8,		// seven segements
	VGA_CLK,   														//	VGA Clock
	VGA_HS,															//	VGA H_SYNC
	VGA_VS,															//	VGA V_SYNC
	VGA_BLANK,														//	VGA BLANK
	VGA_SYNC,														//	VGA SYNC
	VGA_R,   														//	VGA Red[9:0]
	VGA_G,	 														//	VGA Green[9:0]
	VGA_B,															//	VGA Blue[9:0]
	CLOCK_50,                                          // 50 MHz clock
	up,down,left,right, reset, debug, isCollide1, randomNumOut);  

	wire [739 : 0] snake_data;

	output [31:0] debug;
	output isCollide1;
	assign isCollide1 = snake_data[424];
		
	////////////////////////	VGA	////////////////////////////
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK;				//	VGA BLANK
	output			VGA_SYNC;				//	VGA SYNC
	output	[7:0]	VGA_R;   				//	VGA Red[9:0]
	output	[7:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[7:0]	VGA_B;   				//	VGA Blue[9:0]
	input				CLOCK_50;
	input up,down,left,right, reset;

	////////////////////////	PS2	////////////////////////////
	input 			resetn;
	inout 			ps2_data, ps2_clock;
	
	////////////////////////	LCD and Seven Segment	////////////////////////////
	output 			   lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon;
	output 	[7:0] 	leds, lcd_data;
	output 	[6:0] 	seg1, seg2, seg3, seg4, seg5, seg6, seg7, seg8;
	output 	[31:0] 	debug_data_in;
	output   [11:0]   debug_addr;
	
	
	wire [31:0] randomNum;
	output [31:0] randomNumOut;
	assign randomNumOut = randomNum;
	
	
	wire			 clock;
	wire			 lcd_write_en;
	wire 	[31:0] lcd_write_data;
	wire	[7:0]	 ps2_key_data;
	wire			 ps2_key_pressed;
	wire	[7:0]	 ps2_out;	
	
	// clock divider (by 5, i.e., 10 MHz)
	pll div(CLOCK_50,inclock);
	assign clock = CLOCK_50;
	
	// UNCOMMENT FOLLOWING LINE AND COMMENT ABOVE LINE TO RUN AT 50 MHz
	//assign clock = inclock;
	
	// your processor
	//processor myprocessor(clock, ~resetn, /*ps2_key_pressed, ps2_out, lcd_write_en, lcd_write_data,*/ debug_data_in, debug_addr);
	
	
	// keyboard controller
	PS2_Interface myps2(clock, resetn, ps2_clock, ps2_data, ps2_key_data, ps2_key_pressed, ps2_out);
	
	// lcd controller
	lcd mylcd(clock, ~resetn, 1'b1, ps2_out, lcd_data, lcd_rw, lcd_en, lcd_rs, lcd_on, lcd_blon);
	
	// example for sending ps2 data to the first two seven segment displays
	Hexadecimal_To_Seven_Segment hex1(ps2_out[3:0], seg1);
	Hexadecimal_To_Seven_Segment hex2(ps2_out[7:4], seg2);
	
	// the other seven segment displays are currently set to 0
	Hexadecimal_To_Seven_Segment hex3(4'b0, seg3);
	Hexadecimal_To_Seven_Segment hex4(4'b0, seg4);
	Hexadecimal_To_Seven_Segment hex5(4'b0, seg5);
	Hexadecimal_To_Seven_Segment hex6(4'b0, seg6);
	Hexadecimal_To_Seven_Segment hex7(4'b0, seg7);
	Hexadecimal_To_Seven_Segment hex8(4'b0, seg8);
	
	// some LEDs that you could use for debugging if you wanted
	assign leds = 8'b00101011;
	
		
	// VGA
	//wire [1600:0] board;
	//wire [200:0] snake1, snake2;
	//wire head1, head2;
	//wire length1, length2;
	//wire score1, score2;
	//wire stage;
	//wire isDrawing;
	
	//wire [11:0] address_dmem_fromVGA;
	//wire [31:0] data_fromVGA;
	//wire wren_fromVGA;
	//wire [31:0] q_dmem_toVGA;
	
	integer move1, move2, counter;
	reg loadSeed;
	
	initial begin
		move1 = 32'd2;
		move2 = 32'd2;
		counter = 32'd0;
		loadSeed = 1'b1;
	end
	
	
	always@(*) begin
		if (up==1'b0 && move1 != 3) begin
			move1 = 1;
		end
		else if (right==1'b0 && move1 != 4) begin
			move1 = 2;
		end
		else if (down==1'b0 && move1 != 1) begin
			move1 = 3;
		end
		else if (left==1'b0 && move1 != 2) begin
			move1 = 4;
		end
	end
	
	always@(posedge clock) begin
	
		if (counter == 1) begin
			loadSeed = 1'b0;
		end
		counter = counter + 1;
	
	end
	
	
	Reset_Delay			r0	(.iCLK(CLOCK_50),.oRESET(DLY_RST)	);
	VGA_Audio_PLL 		p1	(.areset(~DLY_RST),.inclk0(CLOCK_50),.c0(VGA_CTRL_CLK),.c1(AUD_CTRL_CLK),.c2(VGA_CLK)	);

	
	//snake2 s2 (.clock(VGA_CLK), .rstage(stage), .isDrawing(isDrawing));
	vga_controller vga_ins(.iRST_n(DLY_RST),
								 .iVGA_CLK(VGA_CLK),
								 .oBLANK_n(VGA_BLANK),
								 .oHS(VGA_HS),
								 .oVS(VGA_VS),
								 .b_data(VGA_B),
								 .g_data(VGA_G),
								 .r_data(VGA_R), .up(up), .down(down), .left(left), .right(right),
								 .snake_data(snake_data));
								 //.board(board), 
								 //.snake1(snake1), .snake2(snake2), 
								 //.head1(head1), .head2(head2),
								 //.length1(length1), .length2(length2),
								 //.score1(score1), .score2(score2),
								 //.stage(stage), 
								 //.isDrawing(isDrawing));
								 
	
	 /** IMEM **/
    wire [11:0] address_imem;
    wire [31:0] q_imem;
    imem my_imem(
        .address    (address_imem),            // address of data
        .clock      (~clock),                  // you may need to invert the clock
        .q          (q_imem)                   // the raw instruction
    );

    /** DMEM **/
    wire [11:0] address_dmem;
    wire [31:0] data;
    wire wren;
    wire [31:0] q_dmem;
    dmem my_dmem(
        .address    (/* 12-bit wire */address_dmem),       // address of data
        .clock      (~clock),                  // may need to invert the clock
        .data	    (/* 32-bit data in */data),    // data you want to write
        .wren	    (/* 1-bit signal */wren),      // write enable
        .q          (/* 32-bit data out */q_dmem)    // data from dmem
    );
	 

	 linear_rng lr1 (.clock(clock), .initialSeed(32'b0), .random(randomNum));
	 //rng rng1(.clk(VGA_CLK), .reset(1'b1), .loadseed_i(loadSeed), .rngOut(randomNum[11:0]));
	 //assign randomNum[31:12] = 20'b0;
//	 assign randomNum = 32'b0;
	 
	 
	 /** REGFILE **/
    // Instantiate your regfile
    wire ctrl_writeEnable;
    wire [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
    wire [31:0] data_writeReg;
    wire [31:0] data_readRegA, data_readRegB;
    regfile my_regfile(
        clock,
        ctrl_writeEnable,
        reset,
        ctrl_writeReg,
        ctrl_readRegA,
        ctrl_readRegB,
        data_writeReg,
        data_readRegA,
        data_readRegB,
		  move1, debug, randomNum
    );
	 
	 
	 /** PROCESSOR **/
    processor my_processor(
        // Control signals
        clock,                          // I: The master clock
        reset,                          // I: A reset signal

        // Imem
        address_imem,                   // O: The address of the data to get from imem
        q_imem,                         // I: The data from imem

        // Dmem
        address_dmem,                   // O: The address of the data to get or put from/to dmem
        data,                           // O: The data to write to dmem
        wren,                           // O: Write enable for dmem
        q_dmem,                         // I: The data from dmem

        // Regfile
        ctrl_writeEnable,               // O: Write enable for regfile
        ctrl_writeReg,                  // O: Register to write to in regfile
        ctrl_readRegA,                  // O: Register to read from port A of regfile
        ctrl_readRegB,                  // O: Register to read from port B of regfile
        data_writeReg,                  // O: Data to write to for regfile
        data_readRegA,                  // I: Data from port A of regfile
        data_readRegB,                   // I: Data from port B of regfile
		  snake_data
    );


			
	/*
	snake snake1 (.rboard(board), .clock(VGA_CLK), .reset(reset),
		.rsnake1(snake1), .rsnake2(snake2),
		.rhead1(head1), .rhead2(head2),
		.rlength1(length1), .rlength2(length2),
		.rscore1(score1), .rscore2(score2),
		.rstage(stage),
		.move1(move1), .move2(move2),
		.isDrawing(isDrawing));*/
	
	
endmodule
