	component equal1 is
		port (
			source : out std_logic_vector(0 downto 0);                     -- source
			probe  : in  std_logic_vector(49 downto 0) := (others => 'X')  -- probe
		);
	end component equal1;

	u0 : component equal1
		port map (
			source => CONNECTED_TO_source, -- sources.source
			probe  => CONNECTED_TO_probe   --  probes.probe
		);

